module Mpu (

);

endmodule