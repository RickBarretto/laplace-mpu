module Fetch(
    transmiter, // PIN_E9
    receiver,   // PIN_D9
    RTS,        // PIN_B8
    CTS         // PIN_C8
);


endmodule